
`timescale 1ns/1ps
module arbiter(_req, _frame, _IRDY, clk, _reset,  final_gnt);
input _frame, _IRDY, clk, _reset;
input[2:0] _req;
output[2:0] final_gnt;
integer counter = 0;
reg[2:0] final_gnt, _gnt, req_shifted;
reg[1:0] pointer;
reg currState;

parameter
    IDLE = 1'b0,
    INUSE = 1'b1;
    
    
//---Mini-State Machine--//
//This section was to designed for our state machine. Ideally we simplified our FSM to only have two states, IDLE and INUSE(busy). Because the state of the FSM
//also depended on signals such as Frame#,IRDY#, and RESET#; we included such test cases that would affect the state of the bus. For instance, our State machine 
//takes into account, the case where the requestor is granted the bus, but the requestor has yet to assert its FRAME# signal. A timer(counter) will begin, and
//if Frame# is not asserted within 16 clock cycles, the bus will return to the idle state and the grant vector will reset to not active. Other test cases, include
//when FRAME# and IRDY# are deasserted, the bus will return to the IDLE state, and arbiter can grant another requestor the bus. etc.
always @ (posedge clk, negedge _reset)
begin
//#RESET signal initializes the state of the FSM, priority pointer , and tri-states the request vector.
    if(_reset == 1'b0 )
    begin
        pointer = 0;
        final_gnt = 3'b111;
        req_shifted = 3'bZZZ;
        currState = IDLE;
    end
//Rotate the request vector in order to have the pointed request signal be on the highest priority position. I.E. if 
//the highest priority device pointer is set to Device 1 and the request vector is 101. Then we will need to right shift
// the vector until Bit1 (Device1) is on the highest priority position(0). So the the result will be 110.
     case (pointer)
        2'b00: 
            req_shifted = _req;
        2'b01:
            req_shifted = {_req[0], _req[2:1]};
        2'b10:
            req_shifted = {_req[1:0], _req[2]};
    endcase
//End of Request Signal Rotation//

//----------------------------------Simple Priority Arbiter--------------------------------------------//
//In a simple priority arbiter, each requester is assigned a fixed priority, and the grant is given 
//to the active requester with the highest priority. For example, if the request vector into the arbiter 
//is req[N-1:0], req[0] is typically declared the highest priority. If req[0] is active, it gets the grant.
// If not, and req[1] is active, grant[1] is asserted, and so on. In our design we feed in the shifted/rotated request 
//signal and the arbiter will generate a grant signal. In this example, since the rotated request signal was 110; Our 
// output grant signal from the arbiter should be 110.
	casez (req_shifted)
		3'b??0:
			_gnt = 3'b110;
		3'b?01:
			_gnt = 3'b101;
		3'b011:
			_gnt = 3'b011;

	endcase
//------------------------------------End of Simple Priority Arbiter------------------------------------------//

//Unrotating the grant signal in order to get the final grant request that the arbiter will generate. In order to determine
//the final grant signal, we must "unrotate" the grant  signal that was produced fromt the simple priority arbiter, to grant
// the proper device the bus.
//We must also check the the bus is currently not in use i.e. IDLE, and if it is idle, grant that the requester the bus while also updating
//the priority pointer. 
//In our example, the pointer was still pointing at Device0, so since bit0 is already set at the highest priority, we will not need to unrotate the 
//grant signal generated, and we will only need to set the final grant signal equal to the grant signal generated by the simple priority arbiter. I.E.
//final_gnt = _gnt; and update the pointer to point to Device1 as the device with the highest priority.
 	if(currState == IDLE)
    begin
        case (pointer)
            2'b00:     
              final_gnt = _gnt;
            2'b01:
               final_gnt = { _gnt[1:0], _gnt[2]};
            2'b10:
               final_gnt = {_gnt[0], _gnt[2:1]};
        endcase 
   	end
//------------------------------------End of UnRotating  Request Signal ------------------------------------------//

    //Test case if either FRAME# and IRDY# are deasserted, or timer is over 16 clock cycles, 
    //The current State of the bus will return to idle and the grant signal will reset to not active.
    if((_frame == 1'b1 && _IRDY == 1'b1) || counter > 16)
    begin
        currState = IDLE;
        final_gnt = 3'b111;
        if(counter > 16)
           if(pointer == 2)
        	pointer = 0;
        else 
        	pointer = pointer + 1;
        counter = 0;
    end
    //If frame has not been asserted after grant signal was generated, start the timer. 
    else if(_frame == 1'b1 && final_gnt > 0)
        counter = counter +1;
    //Valdition of Transaction case, once grant signal was outputted, the current State of the bus must be 
    //updated to busy(INUSE).
    else if(currState != INUSE && _frame == 1'b0)
    begin
        currState = INUSE;
        if(pointer == 2)
        	pointer = 0;
        else 
        	pointer = pointer + 1;
        counter = 0;
    end
    //Start timer for Data phase transfer, after address phase has been validated. 
    if(currState == INUSE && counter <= 8)
        counter = counter +1;
    //If transaction is not completed within 8 clock cycles after entering data phase, bus will return to idle state.
    else if(currState == INUSE && counter > 8)
    begin
        currState = IDLE;        
        final_gnt = 3'b111;
    end
    //--------------------------------------------------------END of UnRotating Grant Signal------------------------------------------------------------//
end
//-----------------------------------------------------MONITOR SIGNALS AND DISPLAY DATA----------------------------------------------------------------------//
always @ (posedge clk)
begin
 $timeformat(-9, 0, " ns", 5);
 $display("Current Time: %t\nThe Device with the NEW highest priority is Device%d.\nThe requests signal was:%3b\t_frame: %b\t_IRDY: %b\n",$time, pointer, _req,_frame, _IRDY );
 $display("Current Time: %t\nThe current state of the bus is %b (0 = IDLE, 1 = BUSY)\nThe grant signal was: %3b\n",$time, currState, final_gnt);
//Delay to print the Bus state after monitor Strings have been printed. 
#0.2;
    if(_frame == 1'b1 && _IRDY == 1'b1)
        $display("Current Time:%t\nBus Idle.\n\n",$time);
     else if (_frame == 1'b1 && _IRDY == 1'b0)
        $display("Current Time:%t\nInitiator is ready to complete last data transfer of transaction.But has not been completed.\n\n",$time);
     else if (_frame == 1'b0 && _IRDY == 1'b1)
        $display("Current Time:%t\nA transaction is in progress and the initiator is not ready to complete the current data transfer.\n\n",$time);   
     else if (_frame == 1'b0 && _IRDY == 1'b0)
        $display("Current Time:%t\nA transaction is currently in progress and the initiator is ready to complete it.\n\n",$time);
     else
        $display("Current Time:%t\nBus Idle.\n\n",$time);
end
endmodule